`define Verilator



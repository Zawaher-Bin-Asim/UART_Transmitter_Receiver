`define Vivado

